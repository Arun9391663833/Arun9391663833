module router_reg(clock,resetn,pkt_valid,data_in,fifo_full,rst_int_reg,detect_add,ld_state,laf_state,full_state,lfd_state,parity_done,low_pkt_valid,err,dout);
input clock,resetn,pkt_valid,fifo_full,rst_int_reg,detect_add,ld_state,laf_state,full_state,lfd_state;
input [7:0]data_in;
output reg [7:0]dout;
output reg err,parity_done,low_pkt_valid;
reg [7:0]header,internal_parity,full_state_byte,packet_parity;
//dout logic
always@(posedge clock)
begin
    if(!resetn)
	begin 
	    dout<=8'b0;
	end
	else 
	begin
	    if(detect_add&&pkt_valid&&data_in[1:0]!=3)
		    dout<=dout;
		else
		    if(lfd_state)
			    dout<=header;
			else if(ld_state&&~fifo_full)
			    dout<=data_in;
			else if(ld_state&&fifo_full)
			    dout<=dout;
			else if(laf_state)
			    dout<=full_state_byte;
			else 
			    dout<=dout;
	end
end

//fifo_full_byte
always@(posedge clock)
begin
  if(!resetn)
    full_state_byte<=0;
  else 
  begin
     if(ld_state && fifo_full)
          full_state_byte<=data_in;
      else
         full_state_byte<=full_state_byte;
  end
end

//Header
always@(posedge clock)
begin
  if(!resetn)
    header<=0;
  else 
  begin
    if(detect_add && pkt_valid && (data_in[1:0]!=3))
        header<=data_in;
    else
        header<=header;
  end
end

//parity
always@(posedge clock)
begin
  if(!resetn)
     internal_parity<=0;
  else 
  begin
  if(detect_add)
      internal_parity<=0;
  else if(lfd_state)
      internal_parity<= internal_parity ^ header ;
  else
    if(ld_state && pkt_valid && ~full_state)
        internal_parity<= internal_parity ^data_in;
  end
end

//low_packet_valid
always@(posedge clock)
begin
  if(!resetn)
    low_pkt_valid<=0;
  else 
  begin
    if(rst_int_reg)
        low_pkt_valid<=1'b0;
    else if(ld_state && ~(pkt_valid))
        low_pkt_valid<=1'b1;
    else 
        low_pkt_valid <= low_pkt_valid;
  end
end


//paritydone
always@(posedge clock)
begin
  if(!resetn)
    parity_done<=0;
  else
  begin
    if(detect_add)
    parity_done <= 0;
    else if( (ld_state && ~(pkt_valid) && ~fifo_full) || (laf_state && (low_pkt_valid) && ~parity_done))
          parity_done<=1'b1;
    else
          parity_done<=parity_done;
  end
end

//packet parity
always@(posedge clock)
begin
  if(!resetn)
    packet_parity<=0;
  else if(ld_state && ~pkt_valid)
    packet_parity<=data_in;
  else
    packet_parity<=packet_parity;
end

//error          
always@(posedge clock)
begin
  if(~resetn)
    err <= 0;
  else
    begin  
      if(parity_done)
      begin
        if(internal_parity==packet_parity)
         err<=1'b0;
        else
          err<=1'b1;         
      end
      else
        err<=1'b0;
    end
end

endmodule
